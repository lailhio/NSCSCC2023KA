module datapath(

	input wire clk,rst,
	
	input wire  [5 :0] ext_int, //中断
    
    //inst
    output wire [31:0] PC_IF1,  //Inst addr
    output wire        inst_enF, 
    input wire  [31:0] instr1_F2,  instr2_F2, 
    input wire         i_cache_stall,

    //data
    output wire mem_enE,                    
    output wire [31:0] virtual_data_addrE,     // Write Address
    input  wire [31:0] mem_rdataM,    // Read Data
    output wire [3 :0] mem_write_selectE,      // Write Enable
    output wire [31:0] writedataE,    // Write Data
    input wire         d_cache_stall,
    output wire [1:0] data_size,

    output wire        icache_Ctl, dcache_ctl, 
	//debug interface
    output wire[31:0] debug_wb_pc,
    output wire[3:0] debug_wb_rf_wen,
    output wire[4:0] debug_wb_rf_wnum,
    output wire[31:0] debug_wb_rf_wdata,
    output wire [31:0] debug_cp0_count,
    output wire [31:0] debug_cp0_random,
    output wire [31:0] debug_cp0_cause,
    output wire debug_int,
    output wire debug_commit
    );
	
	//--------InstFetch1 stage----------
	wire [31:0] Pc1Plus4F, Pc1Plus8F, PcPlus12F;    //pc
    wire [31:0] Pc2Plus4F, Pc2Plus8F;
    wire [31:0] PcFlopF;
    
    wire pcErrorF;  // pc错误

    //--------InstFetch2 stage----------
	wire [31:0] Pc1Plus4F2, Pc1Plus8F2, PcPlus12F2;    //pc
    wire [31:0] Pc2Plus4F2, Pc2Plus8F2;
    wire [31:0] PcF2, PcOriF2;    //pc
    wire        delayslot_masterF2, delayslot_slaveF2; // 此时的D阶段（即上一条指令）是否为跳转指令
    wire pcErrorF2;
    wire        branch1F2, jump1F2;
    wire [2:0]  branch_judge_control1F2;
	//----------decode stage---------
    wire pcErrorD;
    ctrl_sign   dec_sign1D, dec_sign2D;
    wire        master_only_oneD, slave_only_oneD;
    wire        master_mem_conflitD, slave_mem_conflitD;
	wire [31:0] instr1D, instr2D;  //指令
    wire [31:0] PcD, PcOriD, Pc1Plus4D, Pc1Plus8D, PcPlus12D;  //pc
    wire [31:0] Pc2Plus4D, Pc2Plus8D;
    wire [31:0] src1_a1D, src1_b1D,src1_aD, src1_bD; //alu输入（操作数
    wire [31:0] src2_a1D, src2_b1D,src2_aD, src2_bD; //alu输入（操作数
    wire [31:0] Mrd1D, Mrd2D, immd1D, pc_branch1D, pc_jump1D;  //寄存器读出数据 立即数 pc分支 跳转
    wire [31:0] Srd1D, Srd2D, immd2D, pc_branch2D, pc_jump2D;  //寄存器读出数据 立即数 pc分支 跳转
    wire        pred_take1D, pred_take2D, branch1D, branch2D, jump1D, jump2D;  //立即数扩展 分支预测 branch jump信号

    wire        delayslot_masterD, delayslot_slaveD;//指令是否在延迟槽
    wire [2:0]  forward1_1D, forward2_1D;
    wire [2:0]  forward1_2D, forward2_2D;
	//-------execute stage----------
    wire pcErrorE;
    ctrl_sign   dec_sign1E, dec_sign2E;
	wire [31:0] PcE, PcOriE, Pc1Plus4E, Pc1Plus8E, PcPlus12E; //pc pc+4 寄存器号 写内存 立即数
    wire [31:0] Pc2Plus4E, Pc2Plus8E;

    wire [31:0] src1_a1E, src1_b1E;
    wire [31:0] src2_a1E, src2_b1E;
    wire [31:0] src1_aE, src1_bE;
    wire [31:0] src2_aE, src2_bE;
    wire [31:0] aluout1E, aluout2E; //alu输出
    wire        branch1E, branch2E; //分支信号
    wire [31:0] pc_branch1E, pc_branch2E;  //分支跳转pc
    wire        pred_failedE, pred_failed_masterE, pred_failed_slaveE;  //分支预测失败
    wire        pred_take1E, pred_take2E;  //分支预测

    wire [31:0] instr1E, instr2E;
    wire        alu_stallE;  //alu暂停
    wire        actual_take1E, actual_take2E;  //分支预测 实际结果
 // 异常处理信号
    wire        addrErrorLw1E, addrErrorLw2E, addrErrorSw1E, addrErrorSw2E; //访存指令异常
    wire        overflow1E, overflow2E; //溢出
    wire        trap1E ,trap2E; //自陷
	
	// cp0	
    wire [31:0] except_type1E, except_type2E;  // 异常类型
    wire        flush_exception_masterE, flush_exception_slaveE;  // 发生异常时需要刷新流水线
    wire [31:0] pc_exception1E, pc_exception2E; //异常处理的地址0xbfc0_0380，若为eret指令 则为返回地址
    wire        pc_trap1E, pc_trap2E; // 发生异常时pc特殊处理
    wire [31:0] badvaddr1E, badvaddr2E;
    wire [31:0] cp0_statusE, cp0_causeE, cp0_epcE, cp0_out1E, cp0_out2E;
	//----------mem stage--------
    wire pcErrorM;
    ctrl_sign   dec_sign1M, dec_sign2M;
	wire [31:0] pcM, PcOriM, Pc2Plus4M;  // pc
    wire [31:0] aluout1M, aluout2M; //alu输出
    wire [31:0] instr1M, instr2M;  //指令
    wire [31:0] result_rdataM;  
    wire [31:0] data_srcM;  
    wire [31:0] result1M, result2M;  // mem out
    wire [31:0] pc_branch1M, pc_branch2M; //分支跳转地址
    wire [31:0] src1_b1M, src2_b1M;
    //异常处理信号 exception
    wire        overflow1M, overflow2M;  //算数溢出
    wire        trap1M, trap2M;  //自陷指令
    wire        addrErrorLw1M, addrErrorLw2M, addrErrorSw1M, addrErrorSw2M; //访存指令异常
    wire        pcErrorM;  //pc异常

	//------writeback stage----------
    wire pcErrorW;
    ctrl_sign   dec_sign1W, dec_sign2W;
	wire [31:0] result1W, result2W;
    wire [31:0] pcW, Pc2Plus4W;
	wire [31:0] instr1W, instr2W;
    
    //------stall sign---------------
    wire stallF, stallF2, stall_masterD, stall_masterE, stall_masterM, stall_masterW ,stallDblank;
    wire stall_slaveD, stall_slaveE, stall_slaveM, stall_slaveW;

    wire flushF, flushF2, flush_masterD, flush_masterE, flush_masterM, flush_masterW;
    wire flush_slaveD, flush_slaveE, flush_slaveM, flush_slaveW, fulsh_ex;
//------------------------------------------Data------------------------------------------
	//--------------------debug---------------------
    assign debug_wb_pc          = (clk) ? pcW : Pc2Plus4W;
    assign debug_wb_rf_wen      = (rst) ? 4'b0000 : ((clk) ? {4{dec_sign1W.regwrite & ~stall_masterW}}: {4{dec_sign2W.regwrite & ~stall_slaveW}});
    assign debug_wb_rf_wnum     = (clk) ? dec_sign1W.writereg : dec_sign2W.writereg;
    assign debug_wb_rf_wdata    = (clk) ? result1W : result2W;
//------------------------------------------Hazard-------------------------------------------
//hazard detection
	hazard hazard0(
        .i_cache_stall(i_cache_stall),
        .d_cache_stall(d_cache_stall),
        .alu_stallE(alu_stallE),
        .master_only_oneD(master_only_oneD), .slave_only_oneD(slave_only_oneD), 
        .master_mem_conflitD(master_mem_conflitD), .slave_mem_conflitD(slave_mem_conflitD),

        .jump1D (jump1D), .jump2D (jump2D), 
        .pred_failed_masterE(pred_failed_masterE), .pred_failed_slaveE(pred_failed_slaveE),
        .flush_exception_masterE(flush_exception_masterE), .flush_exception_slaveE(flush_exception_slaveE),
        .fulsh_ex(fulsh_ex), .Blank1_SL(Blank1_SL), .Blank2_SL(Blank2_SL),

        .dec_sign1D(dec_sign1D), .dec_sign2D(dec_sign2D), 
        .dec_sign1E(dec_sign1E), .dec_sign2E(dec_sign2E), 
        .dec_sign1M(dec_sign1M), .dec_sign2M(dec_sign2M), 
        .dec_sign1W(dec_sign1W), .dec_sign2W(dec_sign2W), 
        .pred_take1D(pred_take1D), .pred_take2D(pred_take2D),

        .rs1D(instr1D[25:21]), .rt1D(instr1D[20:16]),
        .rs2D(instr2D[25:21]), .rt2D(instr2D[20:16]),
        
        // Master
        .stallF(stallF), .stallF2(stallF2), .stall_masterD(stall_masterD), .stall_masterE(stall_masterE), 
        .stall_masterM(stall_masterM), .stall_masterW(stall_masterW),
        // Slave
        .stall_slaveD(stall_slaveD), .stall_slaveE(stall_slaveE), 
        .stall_slaveM(stall_slaveM), .stall_slaveW(stall_slaveW),
        
        // Master
        .flushF(flushF), .flushF2(flushF2), .flush_masterD(flush_masterD), .flush_masterE(flush_masterE), 
        .flush_masterM(flush_masterM), .flush_masterW(flush_masterW),
        // Slave
        .flush_slaveD(flush_slaveD), .flush_slaveE(flush_slaveE), .flush_slaveM(flush_slaveM), 
        .flush_slaveW(flush_slaveW),

        // ctrl
        .stallDblank(stallDblank), .icache_Ctl(icache_Ctl),   .dcache_ctl(dcache_ctl),
        .forward1_1D(forward1_1D), .forward1_2D(forward1_2D), .forward2_1D(forward2_1D), .forward2_2D(forward2_2D)
    );

    //--------------------------------------Fetch------------------------------------------------
    
    assign inst_enF = ~(fulsh_ex) & ~pcErrorF & ~pred_failedE ;
    // pc+4
    assign PcFlopF = {PC_IF1[31:3], 3'b0};
    assign Pc1Plus4F = PcFlopF + 4;
    assign Pc1Plus8F = PcFlopF + 8;
    assign Pc2Plus4F = PcFlopF + 4;
    assign Pc2Plus8F = PcFlopF + 8;
    assign PcPlus12F = PcFlopF + 12;
    assign pcErrorF = |(PC_IF1[1:0] ^ 2'b0) ? 1'b1 : 1'b0; // Whatever Flush all
    // pc reg
    pc_reg pc(
        .clk(clk), .rst(rst), .stallF(stallF),
        .actual_take1E(actual_take1E), .actual_take2E(actual_take2E), .pred_take1E(pred_take1E), .pred_take2E(pred_take2E),
        .pred_take1D(pred_take1D), .pred_take2D(pred_take2D), .pc_trap1E(pc_trap1E),  .pc_trap2E(pc_trap2E), 
        .jump1D(jump1D), .jump2D(jump2D),

        .pc_exception1E(pc_exception1E), .pc_exception2E(pc_exception2E),
        .pc_branch1E(pc_branch1E), .pc_branch2E(pc_branch2E),
        .pc_jump1D(pc_jump1D), .pc_branch1D(pc_branch1D), .pc_jump2D(pc_jump2D), .pc_branch2D(pc_branch2D), 
        .PcPlus8F(Pc1Plus8F), .PcPlus8E(Pc1Plus8E), .PcPlus12E(PcPlus12E), 

        .pc(PC_IF1)
    );
    
	//----------------------------------------InstFetch2------------------------------------------------
    wire inst_enF2;
    wire [31:0] instr1_validF2, instr2_validF2;
    flopstrc #(32) flopPcF2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(PcFlopF),.out(PcF2));
    flopstrc #(32) flopPcOriF2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(PC_IF1),.out(PcOriF2));
    flopstrc #(32) flopPc1Plus4F2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(Pc1Plus4F),.out(Pc1Plus4F2));
    flopstrc #(32) flopPc1Plus8F2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(Pc1Plus8F),.out(Pc1Plus8F2));
    flopstrc #(32) flopPc2Plus4F2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(Pc2Plus4F),.out(Pc2Plus4F2));
    flopstrc #(32) flopPc2Plus8F2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(Pc2Plus8F),.out(Pc2Plus8F2));
    flopstrc #(32) flopPcplus12F2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in(PcPlus12F),.out(PcPlus12F2));
    flopstrc #(2) flopInstEnF2(.clk(clk),.rst(rst),.stall(stallF2),.flush(flushF2),.in({inst_enF, pcErrorF}),.out({inst_enF2, pcErrorF2}));
    assign instr1_validF2 = {32{inst_enF2}} & instr1_F2;  // Discard Not Valid
    assign instr2_validF2 = {32{inst_enF2}} & instr2_F2;  // Discard Not Valid
    predec predecode(.instrF2(instr1_validF2), .branchF2(branch1F2), .jumpF2(jump1F2), .branch_judge_control(branch_judge_control1F2));
    assign delayslot_masterF2 = branch2D | jump2D; //通过前一条指令，判断是否是延迟槽
    assign delayslot_slaveF2 =  branch1F2 | jump1F2; //通过前一条指令，判断是否是延迟槽
    //-----------------------InstFetch2Flop------------------------------


	//----------------------------------------Decode------------------------------------------------
    //-----------------------master---------------------------
    flopstrc #(32) flopPcD(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),.in(PcF2),.out(PcD));
    flopstrc #(32) flopPcOriD(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),.in(PcOriF2),.out(PcOriD));
    flopstrc #(32) flopPc1Plus4D(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),.in(Pc1Plus4F2),.out(Pc1Plus4D));
    flopstrc #(32) flopPc1Plus8D(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),.in(Pc1Plus8F2),.out(Pc1Plus8D));
    flopstrc #(32) flopInst1D(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),.in(instr1_validF2),.out(instr1D));
    flopstrc #(2) flopIsdelay1D(.clk(clk),.rst(rst),.stall(stall_masterD),.flush(flush_masterD),
        .in({delayslot_masterF2, pcErrorF2}),.out({delayslot_masterD, pcErrorD}));
    //-----------------------slave---------------------------
    flopstrc #(32) flopPc2Plus4D(.clk(clk),.rst(rst),.stall(stall_slaveD),.flush(flush_slaveD),.in(Pc2Plus4F2),.out(Pc2Plus4D));
    flopstrc #(32) flopPc2Plus8D(.clk(clk),.rst(rst),.stall(stall_slaveD),.flush(flush_slaveD),.in(Pc2Plus8F2),.out(Pc2Plus8D));
    flopstrc #(32) flopPcplus12D(.clk(clk),.rst(rst),.stall(stall_slaveD),.flush(flush_slaveD),.in(PcPlus12F2),.out(PcPlus12D));
    flopstrc #(32) flopInst2D(.clk(clk),.rst(rst),.stall(stall_slaveD),.flush(flush_slaveD),.in(instr2_validF2),.out(instr2D));
    flopstrc #(1) flopIsdelay2D(.clk(clk),.rst(rst),.stall(stall_slaveD),.flush(flush_slaveD),
        .in({delayslot_slaveF2}),.out({delayslot_slaveD}));
    //-----------------------DecodeFlop----------------------------------
	maindec main_dec1(.instrD(instr1D), .instr2D(instr2D), .dec_sign(dec_sign1D), 
                .only_oneD_inst(master_only_oneD), .Mem_conflit(master_mem_conflitD));
	maindec main_dec2(.instrD(instr2D), .instr2D(instr1D), .dec_sign(dec_sign2D), 
                .only_oneD_inst(slave_only_oneD), .Mem_conflit(slave_mem_conflitD));

    //扩展立即数
    signext signex1(dec_sign1D.sign_ex,instr1D[15:0],immd1D);
    signext signex2(dec_sign2D.sign_ex,instr2D[15:0],immd2D);
	//regfile，                             we3                we4
	regfile rf(clk,rst,stall_masterW,dec_sign1W.regwrite, dec_sign2W.regwrite,
            instr1D[25:21], instr1D[20:16], instr2D[25:21], instr2D[20:16],
            dec_sign1W.writereg, dec_sign2W.writereg, result1W, result2W,
            Mrd1D, Mrd2D, Srd1D, Srd2D);
    // 立即数左移2 + pc+4得到分支跳转地址   
    assign dec_sign1D.delayslot = delayslot_masterD;
    assign dec_sign2D.delayslot = delayslot_slaveD;
    assign pc_branch1D = {immd1D[29:0], 2'b00} + Pc1Plus4D; 
    assign pc_branch2D = {immd2D[29:0], 2'b00} + Pc2Plus8D; 
    // Forward 1
    mux8 #(32) mux8_forward1_1D(Mrd1D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, 32'b0,  
                                forward1_1D, src1_a1D);
    mux8 #(32) mux8_forward1_2D(Mrd2D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, 32'b0,  
                                forward1_2D, src1_b1D);
    // Forward 2
    mux8 #(32) mux8_forward2_1D(Srd1D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, 32'b0,  
                                forward2_1D, src2_a1D);
    mux8 #(32) mux8_forward2_2D(Srd2D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, 32'b0,
                                forward2_2D, src2_b1D);
    // Forward 2
    mux8 #(32) mux8_forbranch1D(Mrd1D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, Pc1Plus8D,  
                                (forward1_1D | {3{jump1D | branch1D}}), src1_aD);
    mux8 #(32) mux8_forbranch2D(Srd1D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, PcPlus12D,
                                (forward2_1D | {3{jump2D | branch2D}}), src2_aD);
                                // Forward 1
    mux8 #(32) mux8_forimm1D(Mrd2D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, immd1D,  
                                (forward1_2D | {3{dec_sign1D.is_imm}}), src1_bD);
    mux8 #(32) mux8_forimm2D(Srd2D, result1W, result2W, result1M, result2M, aluout1E, aluout2E, immd2D,  
                                (forward2_2D | {3{dec_sign2D.is_imm}}), src2_bD);
	// BranchPredict
    BranchPredict branch_predict(
        .clk(clk), .rst(rst),
        .flush_masterD(flush_masterD),.stall_masterD(stall_masterD), .flush_slaveD(flush_slaveD), .stall_slaveD(stall_slaveD),
        .instr1D(instr1D), .instr2D(instr2D), .PcF2(PcF2), .PcPlus4F2(Pc2Plus4F2), .PcE(PcE), .PcPlus4E(Pc2Plus4E),
        .branch1E(branch1E), .branch2E(branch2E),  .actual_take1E(actual_take1E), .actual_take2E(actual_take2E),

        .branch1D(branch1D), .branch2D(branch2D),
        .pred_take1D(pred_take1D) ,.pred_take2D(pred_take2D)
    );
    // jump, assign Logic
    jump_control jump_control(
        .instr1D(instr1D), .instr2D(instr2D),
        .PcPlus4D(Pc1Plus4D), .PcPlus8D(Pc2Plus8D),
        .src1_a1D(src1_a1D), .src2_a1D(src2_a1D),

        .jump1D(jump1D), .jump2D(jump2D),
        .pc_jump1D(pc_jump1D), .pc_jump2D(pc_jump2D) 
    );
	//----------------------------------Execute------------------------------------
    //-----------------------master---------------------------
    flopstrc #(32) flopPcE(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(PcD),.out(PcE));
    flopstrc #(32) flopPcOriE(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(PcOriD),.out(PcOriE));
    flopstrc #(32) flopInst1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(instr1D),.out(instr1E));
    flopstrc #(32) flopSrc1a1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(src1_a1D),.out(src1_a1E));
    flopstrc #(32) flopSrc1b1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(src1_b1D),.out(src1_b1E));
    flopstrc #(32) flopSrc1aE(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(src1_aD),.out(src1_aE));
    flopstrc #(32) flopSrc1bE(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(src1_bD),.out(src1_bE));
    flopstrc #(32) flopPc1Plus4E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(Pc1Plus4D),.out(Pc1Plus4E));
    flopstrc #(32) flopPc1Plus8E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(Pc1Plus8D),.out(Pc1Plus8E));
    flopstrc #(32) flopPcbranch1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(pc_branch1D),.out(pc_branch1E));
    flopstrc #(4) flopSign1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),
        .in({branch1D,pred_take1D,delayslot_masterD, pcErrorD}),
        .out({branch1E,pred_take1E,delayslot_masterE, pcErrorE}));
    flopctrl flopctrl1E(.clk(clk),.rst(rst),.stall(stall_masterE),.flush(flush_masterE),.in(dec_sign1D),.out(dec_sign1E));
    //-----------------------slave---------------------------
    flopstrc #(32) flopInst2E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(instr2D),.out(instr2E));
    flopstrc #(32) flopSrc2a1E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(src2_a1D),.out(src2_a1E));
    flopstrc #(32) flopSrc2b1E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(src2_b1D),.out(src2_b1E));
    flopstrc #(32) flopSrc2aE(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(src2_aD),.out(src2_aE));
    flopstrc #(32) flopSrc2bE(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(src2_bD),.out(src2_bE));
    flopstrc #(32) flopPc2Plus4E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(Pc2Plus4D),.out(Pc2Plus4E));
    flopstrc #(32) flopPc2Plus8E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(Pc2Plus8D),.out(Pc2Plus8E));
    flopstrc #(32) flopPcplus12E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(PcPlus12D),.out(PcPlus12E));
    flopstrc #(32) flopPcbranch2E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(pc_branch2D),.out(pc_branch2E));
    flopstrc #(2) flopSign2E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),
        .in({branch2D, pred_take2D}),
        .out({branch2E, pred_take2E}));
    flopctrl flopctrl2E(.clk(clk),.rst(rst),.stall(stall_slaveE),.flush(flush_slaveE),.in(dec_sign2D),.out(dec_sign2E));
    //-----------------------ExFlop---------------------
	//ALU
    alu_top aluitem(
        //input
        .clk(clk),.rst(rst),.flush_slaveE(flush_slaveE),.flush_masterE(flush_masterE),
        .src1_aE(src1_aE), .src1_bE(src1_bE), .src2_aE(src2_aE), .src2_bE(src2_bE),
        .alucontrolE1(dec_sign1E.alucontrol), .alucontrolE2(dec_sign2E.alucontrol), 
        .fulsh_ex(fulsh_ex), .DivMulEn1(dec_sign1E.DivMulEn), .DivMulEn2(dec_sign2E.DivMulEn), 
        .instr1E(instr1E), .instr2E(instr2E),
        //output
        .alustallE(alu_stallE),.overflow1E(overflow1E), .overflow2E(overflow2E),
        .trap1E(trap1E), .trap2E(trap2E),
        .cp0_out1E(cp0_out1E), .cp0_out2E(cp0_out2E),
        .aluoutE1(aluout1E), .aluoutE2(aluout2E)
    );
    
	//在execute阶段得到真实branch跳转情况
    branch_check branch_check1(
        .branch_judge_controlE(dec_sign1E.branch_judge_control),
        .rs_valueE(src1_a1E),
        .rt_valueE(src1_b1E),
        .actual_takeE(actual_take1E)
    );
    branch_check branch_check2(
        .branch_judge_controlE(dec_sign2E.branch_judge_control),
        .rs_valueE(src2_a1E),
        .rt_valueE(src2_b1E),
        .actual_takeE(actual_take2E)
    );
    //分支预测结果
    
    assign pred_failedE = (pred_take1E ^ actual_take1E) | (pred_take2E ^ actual_take2E);
    assign pred_failed_masterE = pred_take1E ^ actual_take1E;
    assign pred_failed_slaveE = pred_take2E ^ actual_take2E;
    // ---------------MemSign------------------------------
    wire [31:0] data_srcE;
    assign mem_enE = (dec_sign1E.mem_read | dec_sign1E.mem_write)& ~flush_exception_masterE 
            | (dec_sign2E.mem_read | dec_sign2E.mem_write)& ~fulsh_ex; //意外刷新时需要
    wire mem_selE = dec_sign1E.mem_read | dec_sign1E.mem_write;
    wire cpu_data_wr_enE = dec_sign1E.mem_write | dec_sign2E.mem_write;
    // Assign Logical
    wire Blank1_SL = (address1E[31:2] == virtual_data_addrM[31:2]) & dec_sign1E.mem_read &  cpu_data_wr_enM;
    wire Blank2_SL = (address2E[31:2] == virtual_data_addrM[31:2]) & dec_sign2E.mem_read &  cpu_data_wr_enM;
    wire [31:0] address1E = src1_aE + src1_bE;
    wire [31:0] address2E = src2_aE + src2_bE;
    mem_control mem_control(
        .clk(clk),          .rst(rst),
        .instr1E(instr1E), .address1E(address1E), 
        .instr2E(instr2E), .address2E(aluout2E), 
        .mem_selE(mem_selE), .Blank1_SL(Blank1_SL), .stallM(stall_masterM), .flushM(flush_masterM),
        
        .data_wdata1E(src1_b1E),.data_wdata2E(src2_b1E),    //原始的wdata
        .rt_valueM(data_srcM),
        .writedataE(writedataE),
        .mem_write_selectE(mem_write_selectE),
        .data_addrE(virtual_data_addrE), .data_srcE(data_srcE),
        .mem_rdataM(mem_rdataM), .data_rdataM(result_rdataM),
        .data_size(data_size),

        .addr_error_sw1(addrErrorSw1E), .addr_error_lw1(addrErrorLw1E),
        .addr_error_sw2(addrErrorSw2E), .addr_error_lw2(addrErrorLw2E)
    );
    //异常处理
    exception exception1(
        .rst(rst),.ext_int(ext_int),
        //异常信号
        .ri(dec_sign1E.ri), .break_exception(dec_sign1E.breaks), .syscall(dec_sign1E.syscall), 
        .overflow(overflow1E), .addrErrorSw(addrErrorSw1E), .addrErrorLw(addrErrorLw1E), 
        .pcError(pcErrorE), .eretE(dec_sign1E.eret), .trap(trap1E),
        //异常寄存器
        .cp0_status(cp0_statusE), .cp0_cause(cp0_causeE), .cp0_epc(cp0_epcE),
        //记录出错地址
        .PcE(PcOriE),.aluoutE(aluout1E),
        //输出异常处理信号
        .except_type(except_type1E),.flush_exception(flush_exception_masterE),
        .pc_exception(pc_exception1E),
        .pc_trap(pc_trap1E),.badvaddrE(badvaddr1E)
    );
    exception exception2(
        .rst(rst),.ext_int(ext_int),
        //异常信号
        .ri(dec_sign2E.ri), .break_exception(dec_sign2E.breaks), .syscall(dec_sign2E.syscall), 
        .overflow(overflow2E), .addrErrorSw(addrErrorSw2E), .addrErrorLw(addrErrorLw2E), 
        .pcError(pcErrorE), .eretE(dec_sign2E.eret), .trap(trap2E),
        //异常寄存器
        .cp0_status(cp0_statusE), .cp0_cause(cp0_causeE), .cp0_epc(cp0_epcE),
        //记录出错地址
        .PcE(PcOriE),.aluoutE(aluout2E),
        //输出异常处理信号
        .except_type(except_type2E),.flush_exception(flush_exception_slaveE),
        .pc_exception(pc_exception2E),
        .pc_trap(pc_trap2E),.badvaddrE(badvaddr2E)
    );
     // cp0 todo 
    cp0_reg cp0(
        .clk(clk) , .rst(rst),
        .stall_masterW(stall_masterW), .we1_i(dec_sign1E.cp0_write) , .we2_i(dec_sign2E.cp0_write) ,
        .waddr1_i(instr1E[15:11]) , .raddr1_i(instr1E[15:11]), .waddr2_i(instr2E[15:11]) , .raddr2_i(instr2E[15:11]),
        .data1_i(src1_b1E), .data2_i(src2_b1E), .int_i(ext_int),
        .excepttype1_i(except_type1E) , .excepttype2_i(except_type2E), 
        .current_inst_addr1_i(PcOriE), .current_inst_addr2_i(Pc2Plus4E),
        .is_in_delayslot1_i(dec_sign1E.delayslot) , .is_in_delayslot2_i(dec_sign2E.delayslot), 
        .bad_addr1_i(badvaddr1E), .bad_addr2_i(badvaddr2E),
        .status_o(cp0_statusE) , .cause_o(cp0_causeE) ,
        .epc_o(cp0_epcE), .data1_o(cp0_out1E), .data2_o(cp0_out2E)
    );
    
	//-------------------------------------Memory----------------------------------------
    wire [31:0] virtual_data_addrM;
    wire        cpu_data_wr_enM;
    //-----------------------master---------------------------
	flopstrc #(32) flopPcM(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(PcE),.out(pcM));
	flopstrc #(32) flopPcOriM(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(PcOriE),.out(PcOriM));
	flopstrc #(32) flopAlu1M(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(aluout1E),.out(aluout1M));
	flopstrc #(32) flopRtvalue1M(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(src1_b1E),.out(src1_b1M));
    flopstrc #(32) flopRtvalueM(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(data_srcE),.out(data_srcM));
	flopstrc #(32) flopInstr1M(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(instr1E),.out(instr1M));
	flopstrc #(32) flopAddrM(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(virtual_data_addrE),.out(virtual_data_addrM));
    flopstrc #(6) flopSign1M(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),
        .in({overflow1E, trap1E, pcErrorE, addrErrorLw1E, addrErrorSw1E, cpu_data_wr_enE}),
        .out({overflow1M, trap1M, pcErrorM, addrErrorLw1M, addrErrorSw1M, cpu_data_wr_enM}));
    flopctrl flopctrl1M(.clk(clk),.rst(rst),.stall(stall_masterM),.flush(flush_masterM),.in(dec_sign1E),.out(dec_sign1M));
    //-----------------------slave---------------------------
	flopstrc #(32) flopPc2Plus4M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),.in(Pc2Plus4E),.out(Pc2Plus4M));
	flopstrc #(32) flopAlu2M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),.in(aluout2E),.out(aluout2M));
	flopstrc #(32) flopRtvalue2M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),.in(src2_b1E),.out(src2_b1M));
	flopstrc #(32) flopInstr2M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),.in(instr2E),.out(instr2M));
    flopstrc #(4) flopSign2M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),
        .in({overflow2E, trap2E, addrErrorLw2E, addrErrorSw2E}),
        .out({overflow2M, trap2M, addrErrorLw2M, addrErrorSw2M}));
    flopctrl flopctrl2M(.clk(clk),.rst(rst),.stall(stall_slaveM),.flush(flush_slaveM),.in(dec_sign2E),.out(dec_sign2M));
    //----------------------MemoryFlop------------------------
    

    //在aluout1W, cp0_outW 中选择写入寄存器的数据 Todo
    mux2 #(32) mux2_memtoreg1M(aluout1M, result_rdataM,dec_sign1M.mem_read, result1M);
    mux2 #(32) mux2_memtoreg2M(aluout2M, result_rdataM,dec_sign2M.mem_read, result2M);
     
	//-------------------------------------Memory2-------------------------------------------------
    // todo M2 flop
    //-----------------------master---------------------------
	flopstrc #(32) flopPc1W(.clk(clk),.rst(rst),.stall(stall_masterW),.flush(flush_masterW),.in(pcM),.out(pcW));
	flopstrc #(32) flopInstr1W(.clk(clk),.rst(rst),.stall(stall_masterW),.flush(flush_masterW),.in(instr1M),.out(instr1W));
	flopstrc #(32) flopRes1W(.clk(clk),.rst(rst),.stall(stall_masterW),.flush(flush_masterW),.in(result1M),.out(result1W));
    flopctrl flopctrl1W(.clk(clk),.rst(rst),.stall(stall_masterW),.flush(flush_masterW),.in(dec_sign1M),.out(dec_sign1W));
    //-----------------------slave---------------------------
	flopstrc #(32) flopRes2W(.clk(clk),.rst(rst),.stall(stall_slaveW),.flush(flush_slaveW),.in(result2M),.out(result2W));
	flopstrc #(32) flopPc2W(.clk(clk),.rst(rst),.stall(stall_slaveW),.flush(flush_slaveW),.in(Pc2Plus4M),.out(Pc2Plus4W));
	flopstrc #(32) flopInstr2W(.clk(clk),.rst(rst),.stall(stall_slaveW),.flush(flush_slaveW),.in(instr2M),.out(instr2W));
    flopctrl flopctrl2W(.clk(clk),.rst(rst),.stall(stall_slaveW),.flush(flush_slaveW),.in(dec_sign2M),.out(dec_sign2W));
	//------------------Memory2_Flop--------------------------
	
endmodule
